module sevevenseg(hex1,hex0,x,y);

input wire [3:0] x,y;
output wire [6:0] hex1,hex0;

assign hex1[6] = (x[3]&x[2])|(x[3]&x[1])|(~x[3]&~x[2]&~x[1])|(x[2]&x[1]&x[0]);
assign hex1[5] = (x[3]&x[2])|(x[3]&x[1])|(~x[3]&~x[2]&x[0])|(~x[2]&x[1]);
assign hex1[4] = (x[3]&x[2])|(x[3]&x[1])|(x[0])|(x[2]&~x[1]);
assign hex1[3] = (x[2]&~x[1]&~x[0])|(x[2]&x[1]&x[0])|(~x[3]&~x[2]&~x[1]&x[0])|(x[3]&x[2])|(x[3]&x[1]);
assign hex1[2] = (x[3]&x[2])|(x[3]&x[1])|(~x[2]&x[1]&~x[0]);
assign hex1[1] = (x[3]&x[2])|(x[3]&x[1])|(x[2]&~x[1]&x[0])|(x[2]&x[1]&~x[0]);
assign hex1[0] = (x[3]&x[2])|(x[3]&x[1])|(~x[3]&~x[2]&~x[1]&x[0])|(x[2]&~x[1]&~x[0]);

assign hex0[6] = (y[3]&y[2])|(y[3]&y[1])|(~y[3]&~y[2]&~y[1])|(y[2]&y[1]&y[0]);
assign hex0[5] = (y[3]&y[2])|(y[3]&y[1])|(~y[3]&~y[2]&y[0])|(~y[2]&y[1]);
assign hex0[4] = (y[3]&y[2])|(y[3]&y[1])|(y[0])|(y[2]&~y[1]);
assign hex0[3] = (y[2]&~y[1]&~y[0])|(y[2]&y[1]&y[0])|(~y[3]&~y[2]&~y[1]&y[0])|(y[3]&y[2])|(y[3]&y[1]);
assign hex0[2] = (y[3]&y[2])|(y[3]&y[1])|(~y[2]&y[1]&~y[0]);
assign hex0[1] = (y[3]&y[2])|(y[3]&y[1])|(y[2]&~y[1]&y[0])|(y[2]&y[1]&~y[0]);
assign hex0[0] = (y[3]&y[2])|(y[3]&y[1])|(~y[3]&~y[2]&~y[1]&y[0])|(y[2]&~y[1]&~y[0]);

endmodule
