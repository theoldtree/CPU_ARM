module REG #(parameter BITWIDTH = 32) (	
	input wire	CLK,
	input wire	RST,
	input wire	EN,
	input wire	[BITWIDTH - 1:0]	D,
	output reg	[BITWIDTH - 1:0]	Q
); // ???? ??(CLK), ??(RST), EN?, ??(D), ?? Q?? ??

	always @ (posedge CLK) // CLK??? ??????
	begin
		if (RST)		Q<=0; // ????? ??? ??? 0
		else if (EN)	Q<=D; // EN??? 1?? ??? ???
	end
endmodule
