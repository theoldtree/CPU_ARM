
module NZCV_REG #(parameter BITWIDTH = 4)(
	input wire CLK,
	input wire RST,
	input wire [3:0] EN,
	input wire [3:0] D,
	output wire [3:0] Q
);// ???? CLK(??), RST(??), 4??? EN(enable), D(???)? ???? ???? Q(???) ??
reg [3:0] d;
wire en;
// ??? ?? ??? d ? D flipflop? ???? en??
assign en = |EN; // en? ? ??
REG #(BITWIDTH) NZCV (
	.CLK (CLK),
	.RST (RST),
	.EN (en),
	.D (d),
	.Q (Q)
); // REG? ???? ??
always @ (EN) 
	case (EN) 
	4'b0000 : d = Q;
	4'b1110 : d = {D[3:1],Q[0]};
	4'b1111 : d = D;
endcase
// EN? ????? ?? ?? d ? ?? ??? ? ??

endmodule
