`timescale 10ns/1ps
module TB_NZCV_REG;
	reg [3:0] D;
	reg [3:0] EN;
	reg CLK;
	reg RST;
	wire [3:0] Q; // ???? ??? ??? ??? ??
	initial CLK = 1'b0;
	always #1 CLK = ~CLK; // ????
NZCV_REG #(4) NZCV_REG(
	.CLK (CLK),
	.RST (RST),
	.EN (EN),
	.D (D),
	.Q (Q)
); // NZCV_REG? ???? ??
initial
begin
	RST = 1'b1; // ?? ??
	#2
	RST = 1'b0;
	#2
	EN=4'b1111;
	D=4'b1010;
	#2
	EN=4'b1110;
	D=4'b0011;
	#2
	EN=4'b0000;
	D=4'b1111;
	// ??? ??? ?? EN??? D??? ???? ?? ??? ????.
	#2
	$finish();
end

endmodule
